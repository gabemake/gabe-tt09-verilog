//typedef enum states { IDLE, COUNTING, SCORE1, SCORE2, SCORE3, SCORE4, SCOREB, OVER1, OVER2, OVER3, OVER4, OVERB} states_t;
parameter IDLE = 'd 0;
parameter COUNTING = 'd 1;
parameter SCORE1 = 'd 2;
parameter SCORE2 = 'd 3;
parameter SCORE3 = 'd 4;
parameter SCORE4 = 'd 5;
parameter SCOREB = 'd 6;
parameter OVER1 = 'd 7;
parameter OVER2 = 'd 8;
parameter OVER3 = 'd 9;
parameter OVER4 = 'd 10;
parameter OVERB = 'd 11;

//typedef enum display {d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, dB, dV, dE, dR, dD} display_t;
parameter d0 = 'd 0;
parameter d1 = 'd 1;
parameter d2 = 'd 2;
parameter d3 = 'd 3;
parameter d4 = 'd 4;
parameter d5 = 'd 5;
parameter d6 = 'd 6;
parameter d7 = 'd 7;
parameter d8 = 'd 8;
parameter d9 = 'd 9;
parameter dB = 'd 10;
parameter dV = 'd 11;
parameter dE = 'd 12;
parameter dR = 'd 13;
parameter dD = 'd 14;
